package alu_pkg;
  `include "defines.sv"          // common definitions if exists
  `include "alu_transaction.sv"  // transaction class
  `include "alu_generator.sv"    // generator class
  `include "alu_driver.sv"       // driver class
  `include "alu_monitor.sv"      // monitor class
  `include "alu_reference.sv"  // reference model
  `include "alu_scoreboard.sv"   // scoreboard for checking
  `include "alu_environments.sv" // test environment
  `include "alu_test.sv"         // test cases
endpackage
